module lock(
 input [3:0] password_in,  //輸入設定密碼
 input [3:0] password_try,  //輸入猜測密碼
 input      set,     //設定密碼
 input      unlock,    //嘗試解鎖
 output [3:0] password_out,  //目前密碼 
 output reg unlock_out,   //解鎖燈號
 output reg  lock_out,   //上鎖燈號
 output reg  beep=0,     //蜂鳴器
 
 output reg [7:0] R_color, G_color, B_color,
 output reg [3:0] column,  //8*8矩陣
 input CLK
 
 );
 reg [3:0] password;     //儲存密碼
 reg [3:0] count;     //計算時間
 reg check=0;       //在try的時候判斷是否正確
 
 assign password_out = password;  //顯示燈號

 
 divfreq F1(CLK, CLK_div);



initial 
 begin 
  unlock_out=0;
  lock_out=0;
  count=4'b0000;
  R_color=8'b11111111;
  G_color=8'b11111111;
  B_color=8'b11111111;
  column=4'b1000;
 end

 
 
always @(set,unlock)
 begin
  if(set && password_try==4'b1010)  //安全碼1010
   begin
    password = password_in;
    lock_out = 1;
    unlock_out = 0;
    check = 0;   //上鎖狀態
    beep =0 ;
   end
	
  else if(unlock)
   begin 
    if(password_try == password)  //輸入正確
     begin
      lock_out = 0;
      unlock_out = 1;
      check = 1;  //解鎖狀態
      beep =0;
     end
    
    else if(password_try != password )  //輸入錯誤
     begin
       lock_out = 1;
       unlock_out = 0;
       check = 0;
       beep =1;  //蜂鳴器響
     end
   end
 end

 

always@(posedge CLK_div)
if(check) //正確
 begin 
  count <= count + 1'b1;
  if(count>4'b1111)
   count<=4'b1000;
  else if(count==4'b1000) 
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1001)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b11011111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1010)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b10110011;
    B_color<=8'b11111111;
   end
  else if(count==4'b1011)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b10111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1100)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b10111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1101)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b10110011;
    B_color<=8'b11111111;
   end
  else if(count==4'b1110)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b11011111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1111)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
 end
 
 
 
else if(~check) //錯誤
 begin 
  count <= count + 1'b1;
  if(count>4'b1111)
   count<=4'b1000;
  else if(count==4'b1000) 
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1001)
   begin
    column<=count;
    R_color<=8'b10111111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1010)
   begin
    column<=count;
    R_color<=8'b11010011;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1011)
   begin
    column<=count;
    R_color<=8'b11011111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1100)
   begin
    column<=count;
    R_color<=8'b11011111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1101)
   begin
    column<=count;
    R_color<=8'b11010011;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1110)
   begin
    column<=count;
    R_color<=8'b10111111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end
  else if(count==4'b1111)
   begin
    column<=count;
    R_color<=8'b11111111;
    G_color<=8'b11111111;
    B_color<=8'b11111111;
   end  
 end

endmodule



module divfreq(input CLK,output reg CLK_div); //除頻器
reg[24:0] Count;
always@(posedge CLK)
 begin
  if(Count > 1000)
   begin
    Count <= 25'b0;
    CLK_div<=~CLK_div;
   end
  else
   Count<=Count+1'b1;
  end
endmodule